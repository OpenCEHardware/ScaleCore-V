package hsv_core_pkg;

endpackage
